module init