module reg_cont

// Import reg_init, so we can initialize registers here.
import init.reg_init

const sigma := reg_init.init_spregisters()